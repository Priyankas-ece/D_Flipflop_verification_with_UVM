//dff UVM tb interface

//Interface creation for signals
interface dff_interface(input logic clk) ; 
  logic rst;
  logic din;
  logic dout;
endinterface